`timescale 1ns / 1ps

module CPU(
    input clk,
    input rst
);

// Internal Wires
wire [31:0] alu_operand;
wire [31:0] alu_otp;
wire [31:0] pc_instaddr;
wire [31:0] instruction;
wire [31:0] sign_extend;
wire [31:0] reg1data;
wire [31:0] reg2data;
wire [31:0] regwrdata;
wire [31:0] data_mem_in;
wire [31:0] data_mem_out;

wire [1:0]  pcControl;
wire [2:0]  alu_op;
wire [4:0]  reg_radd0;
wire [4:0]  reg_radd1;
wire [4:0]  reg_waddr;
wire [5:0]  alu_control_otp;

wire        reg_wr_add_control;
wire        datamem_readen;
wire        datawr_select;
wire        datamemwriteen;
wire        alusrcselect;
wire        reg_wr_en;
wire        branch_control;
wire        jump_control;
wire        alu_zero;
wire        overflow_signal;

// Program Counter
ProgramCounter prcount (
    .clk(clk),
    .reset(rst),
    .zero(alu_zero),
    .branch(branch_control),
    .jump(jump_control),
    .jumpAddress(instruction[25:0]),
    .branchOffset(instruction[15:0]),
    .regAddress(reg1data),
    .pc(pc_instaddr)
);

// Instruction Memory
InstructionMemoryModule instructionMemory (
    .clk(clk),
    .address(pc_instaddr),
    .readEnable(1'b1),
    .writeEnable(1'b0),
    .dataIn(32'h000000),
    .dataOut(instruction)
);

// Control Unit
control_unit signals (
    .instruction(instruction),
    .RegDst(reg_wr_add_control),
    .MemRead(datamem_readen),
    .MemToReg(datawr_select),
    .ALUOp(alu_op),
    .MemWrite(datamemwriteen),
    .ALUSrc(alusrcselect),
    .RegWrite(reg_wr_en),
    .Branch(branch_control),
    .Jump(jump_control)
);

// Register Read Addresses
assign reg_radd0 = instruction[25:21];
assign reg_radd1 = instruction[20:16];

// Register Write Destination Selection
regmux2x1 reg_wr_dst (
    .select(reg_wr_add_control),
    .in0(reg_radd1),
    .in1(instruction[15:11]),
    .out(reg_waddr)
);

// Register File
Register_File regfile (
    .clk(clk),
    .read_addr1(reg_radd0),
    .read_addr2(reg_radd1),
    .write_addr(reg_waddr),
    .write_data(regwrdata),
    .write_enable(reg_wr_en),
    .read_data1(reg1data),
    .read_data2(reg2data)
);

// Sign Extension
signExtension sign (
    .in(instruction[15:0]),
    .out(sign_extend)
);

// ALU Source Selection
mux2x1 alusrc_select (
    .select(alusrcselect),
    .in0(reg2data),
    .in1(sign_extend),
    .out(alu_operand)
);

// ALU Control
alu_control alucntrl (
    .instruction(instruction),
    .ALUOp(alu_op),
    .ALUFn(alu_control_otp)
);

// ALU
ALU alu (
    .clk(clk),
    .a(reg1data),
    .b(alu_operand),
    .alufn(alu_control_otp),
    .otp(alu_otp),
    .zero(alu_zero),
    .overflow(overflow_signal)
);

// Data Memory
MainMemoryModule data_mem (
    .clk(clk),
    .address(alu_otp),
    .readEnable(datamem_readen),
    .writeEnable(datamemwriteen),
    .dataIn(data_mem_in),
    .dataOut(data_mem_out)
);

// Write Data Selection
mux2x1 write_select (
    .select(datawr_select),
    .in1(data_mem_out),
    .in0(alu_otp),
    .out(regwrdata)
);

// Data Memory Input Assignment
assign data_mem_in = reg2data;

// Debugging Display
always @(posedge clk) begin
    $display("reg_radd0 = %d | reg_radd1 = %d", reg_radd0, reg_radd1);
    $display("INSTRUCTION = %h | reg1data = %h | reg2data = %h | alu_control_otp = %d | datamemwriteen = %d | data_mem_in = %d | alu_otp = %h",
        instruction, 
        reg1data, 
        reg2data,
        alu_control_otp,
        datamemwriteen,
        data_mem_in,
        alu_otp
    );
end

endmodule
